module normalizer (
    input [9:0] in,
    input enable,            // ???? 1 ? ??????????? ????????????
    output [9:0] out
);

    assign out = enable ? (in >> 1) : in;

endmodule
